module adder_16b(
input [7:0] a,
input [15:0] b,
output [15:0] sum);

	assign sum = a+b; //Inputs only
	
endmodule


